progress a3s1
player entities/columbiare 893 1120
world world/world.wld
section com.glowingpigeon.columbiare.state.premade.A3
npc stand 6114 464 entities/npcs/amia.npc dead
npc stand 320 64 entities/npcs/fara.npc
npc stand 896 1056 entities/npcs/test.npc
