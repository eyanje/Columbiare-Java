progress a1s1
player entities/columbiare 454 342
world world/world.wld
section com.glowingpigeon.columbiare.state.premade.A1S1_1
npc stand 320 320 entities/npcs/elder.npc
npc stand 1024 0 entities/npcs/fara.npc
npc stand 0 128 entities/npcs/test.npc
npc stand 0 -512 entities/npcs/amia.npc
